//////////////////////////////////////////////////////////////////////////////////
// Engineer: Robert Wu
// 
// Create Date: 05/01/2019 11:24:22 AM
// Project Name: Single Cycle CPU with 31 Instructions Based on MIPS Architecture
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module extend_cut(
    input [31:0] data_in,
    input [2:0] EC_CS,
    input SIGN_EC,
    output [31:0] data_out
    );
    
    reg [31:0] temp;
    
    always @ (*) begin
        case(EC_CS)
            3'b001: temp <= {(SIGN_EC && data_in[15]) ? 16'hffff : 16'h0000, data_in[15:0]};
            3'b010: temp <= {(SIGN_EC && data_in[7]) ? 24'hffffff : 24'h000000, data_in[7:0]};
            3'b011: temp <= {24'h000000, data_in[7:0]};
            3'b100: temp <= {16'h0000, data_in[15:0]};
            default: temp <= data_in;
        endcase
    end
    
    assign data_out = temp;
    
endmodule

